class washing_machine_transaction extends uvm_sequence_item;
