interface washing_machine_if(input bit clk, input bit rst_n);
